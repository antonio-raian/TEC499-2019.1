
module Problema1Qsys (
	botoes_export,
	clk_clk,
	leds_export,
	reset_reset_n);	

	input	[3:0]	botoes_export;
	input		clk_clk;
	output	[4:0]	leds_export;
	input		reset_reset_n;
endmodule
